module top_module();
    wire a, b, c, d;
endmodule
